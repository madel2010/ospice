
V1 n1 0 1
R1 n1 n2 2
L1 n2 n3 1
C1 n2 0 1

.tran 1 1
